module bin2seg (
    input [3:0] bin_data, //Binary input data
    output [7:0] seg_out //7-segment output data (index 7 is don't care)
    );

// **** TODO **** //



// ************** // 

endmodule
