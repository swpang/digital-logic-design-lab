module bcd_counter(
    input clk, // When clk is rising edge, the counter works.
    input rstn, //When rstn is falling edge, the counter resets.
    input i_toggle, //Active low
    output [3:0] data_out //Binary output
    );

// **** TODO **** //



// ************** // 

endmodule